ENTITY NAND_4 IS
PORT(
	A, B : IN BIT;
	Y : OUT BIT
);
END NAND_4;

ARCHITECTURE NAND_INNER OF NAND_4 IS
SIGNAL X1 : BIT;
SIGNAL X2 : BIT;
SIGNAL X3 : BIT;
BEGIN
	X1 <= NOT (A AND B);
	X2 <= NOT (A AND X1);
	X3 <= NOT (B AND X1);
	Y <= NOT (X2 AND X3);
END NAND_INNER;
