ENTITY BC IS
PORT(
	A, B : IN BIT;
	X, Y, Z : OUT BIT
);
END BC;
ARCHITECTURE BC_INNER OF BC IS
BEGIN
	X <= A AND NOT B;
	Y <= NOT (A XOR B);
	Z <= NOT A AND B;
END BC_INNER;
