
LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
ENTITY DECODER_7447 IS
PORT(
	I : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	X : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
);
END DECODER_7447;

ARCHITECTURE DECODER OF DECODER_7447 IS 
	SIGNAL DECODE : STD_LOGIC_VECTOR(6 DOWNTO 0);
	BEGIN
		PROCESS(I)
		BEGIN
			CASE I IS
				WHEN "0000" => DECODE <= "1111110";
				WHEN "0001" => DECODE <= "0110000";
				WHEN "0010" => DECODE <= "1101101";
				WHEN "0011" => DECODE <= "1111001";
				WHEN "0100" => DECODE <= "0110011";
				WHEN "0101" => DECODE <= "1011011";
				WHEN "0110" => DECODE <= "1011111";
				WHEN "0111" => DECODE <= "1110000";
				WHEN "1000" => DECODE <= "1111111";
				WHEN "1001" => DECODE <= "1111011";
				WHEN OTHERS => NULL; 
			END CASE;
		END PROCESS;
	X <= DECODE;
END DECODER;