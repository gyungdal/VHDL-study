LIBRARY  IEEE;
USE  IEEE.STD_LOGIC_1164.ALL;
USE  IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY  TB_COUNT_8BIT IS
END  TB_COUNT_8BIT;
ARCHITECTURE  HB OF TB_COUNT_8BIT IS
COMPONENT COUNT_8BIT
PORT (
     RESETN : IN STD_LOGIC;
     CLK : IN STD_LOGIC;
     COUNT_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;
SIGNAL RESETN : STD_LOGIC := '0';
SIGNAL CLK : STD_LOGIC := '0';
SIGNAL COUNT_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
BEGIN
PROCESS
BEGIN
     WAIT FOR 10 NS;
     CLK <= NOT CLK;
END PROCESS;
RESETN <= '0', '1' AFTER 15NS, '0' AFTER 500NS, '1' AFTER 550NS;
U_COUNT_8BIT : COUNT_8BIT
PORT MAP (
     RESETN => RESETN,
     CLK => CLK,
     COUNT_OUT => COUNT_OUT
);
END HB;