--TB_HB_83ENCODER.VHD 
LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY TB_HB_83ENCODER IS
END TB_HB_83ENCODER; 
ARCHITECTURE HB OF TB_HB_83ENCODER IS
COMPONENT HB_83ENCODER 
PORT (
     A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
     O : OUT STD_LOGIC_VECTOR(2 DOWNTO 0) 
); 
END COMPONENT; 
SIGNAL A : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000"; 
SIGNAL O : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000"; 
BEGIN 
         A <= "10000000", "01000000" AFTER 100NS, "00100000" AFTER 200NS, "00010000" 
                  AFTER 300NS, "00001000" AFTER 400NS, "00000100" AFTER 500NS, "00000010" 
                  AFTER 600NS, "00000001" AFTER 700NS; 
U_HB_83ENCODER : HB_83ENCODER 
PORT MAP (
         A => A, 
         O => O 
); 
END HB; 	
