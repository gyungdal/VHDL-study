LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY TB_7447 IS
END TB_7447; 
ARCHITECTURE HB OF TB_7447 IS
COMPONENT DECODER_7447 
PORT (
     I : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
     X : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) 
); 
END COMPONENT; 
SIGNAL I : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000"; 
SIGNAL X : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000"; 
BEGIN
        I <= "0000", "0001" AFTER 100NS, "0010" AFTER 200NS, "0011" 
                  AFTER 300NS, "0100" AFTER 400NS, "0101" AFTER 500NS, "0110" 
                  AFTER 600NS, "0111" AFTER 700NS, "1000" AFTER 800NS, "1001" AFTER 900NS; 
U_DECODER_7447 : DECODER_7447 
PORT MAP (
         I => I, 
         X => X 
); 
END HB; 	