LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY TB_HB_2MUX IS 
END TB_HB_2MUX; 
ARCHITECTURE HB OF TB_HB_2MUX IS 
COMPONENT HB_2MUX 
PORT ( 
	I0, I1, S : IN STD_LOGIC; 
	Z : OUT STD_LOGIC 
); 
END COMPONENT; 
SIGNAL I0, I1, S : STD_LOGIC := '0'; 
SIGNAL Z : STD_LOGIC := '0'; 	
BEGIN 
PROCESS 
BEGIN 
WAIT FOR 10NS; 
I0 <= NOT I0; 
END PROCESS; 
PROCESS
 BEGIN WAIT FOR 20NS;
 I1 <= NOT I1; 
END PROCESS;
 S <= '0', '1' AFTER 200NS; 
U_HB_2MUX : HB_2MUX PORT MAP ( I0 => I0, I1 => I1, S => S, Z => Z ); 
END HB; 