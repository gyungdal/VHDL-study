--TB_HB_4FA.VHD 
LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY TB_HB_4FA IS 
END TB_HB_4FA; 
ARCHITECTURE HB OF TB_HB_4FA IS 
COMPONENT HB_4FA 
PORT ( 
        CI : IN STD_LOGIC; 
        A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
        S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
        CO : OUT STD_LOGIC 
); 
END COMPONENT; 
SIGNAL CI : STD_LOGIC := '0'; 
SIGNAL A, B : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000"; 
SIGNAL S: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000"; 
SIGNAL CO : STD_LOGIC := '0'; 
BEGIN 
A <= "0000", "1010" AFTER 200NS, "1111" AFTER 400NS; 
B <= "0000", "1011" AFTER 200NS; 
CI <= '0', '1' AFTER 300NS, '0' AFTER 500NS; 
U_HB_4FA : HB_4FA 
PORT MAP ( 
        CI => CI, 
        A => A, 
        B => B, 
        S => S, 
        CO => CO 
); 
END HB; 