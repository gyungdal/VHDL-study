
LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
ENTITY HB_NOR IS
PORT(
	A, B : IN BIT;
	X : OUT BIT
);
END HB_NOR;

ARCHITECTURE HB OF HB_NOR IS
BEGIN
X <= NOT (A OR B);
END HB;