
LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
ENTITY HB_NAND IS
PORT(
	A, B : IN BIT;
	X : OUT BIT
);
END HB_NAND;

ARCHITECTURE HB OF HB_NAND IS
BEGIN
X <= NOT (A AND B);
END HB;