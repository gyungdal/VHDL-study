LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY TB_HB_38DECODER IS 
END TB_HB_38DECODER;
ARCHITECTURE HB OF TB_HB_38DECODER IS
COMPONENT HB_38DECODER 
PORT (
        A, B, C : IN STD_LOGIC; 
        O : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) ); 
END COMPONENT; 
SIGNAL A, B, C : STD_LOGIC := '0'; 
SIGNAL O : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000"; 
BEGIN 
A <= '0', '1' AFTER 800NS; 
B <= '0', '1' AFTER 400NS, '0' AFTER 800NS, '1' AFTER 1200NS; 
C <= '0', '1' AFTER 200NS, '0' AFTER 400NS, '1' AFTER 600NS, '0' AFTER 800NS, '1' AFTER  
         1000NS, '0' AFTER 1200NS, '1' AFTER 1400NS; 
U_HB_38DECODER : HB_38DECODER 
PORT MAP (
      A => A, 
      B => B, 
      C => C, 
      O => O 
);
 END HB;
